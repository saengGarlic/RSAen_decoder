
module MIPS_top();
	
	wire [11:0] ctrl_wire;
	wire 